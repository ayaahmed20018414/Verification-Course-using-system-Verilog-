package Adder_package; 
`include "driver.svh"
`include "monitor_input.svh"
`include "monitor_output.svh"
`include "Check_output.svh"
endpackage 
