package adder_pkg;
`include "transaction.svh"
`include "generator.svh"
`include "driver.svh"
`include "monitor.svh"
`include "scoreboard.svh"
`include "coverpoint.svh"
endpackage
